`define TXNS 3 
`define SLAVES 1

`define ADDR_WIDTH 8

`define DATA_WIDTH 32 

`define PSEL_WIDTH 4






































